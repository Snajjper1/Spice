* Circuit with one DC Voltage source and 3 resistors in series

vsupply 1 0 dc 22;
r1 2 1 5k;
r2 3 2 3.3k;
r3 3 0 1.2k;

.dc vsupply 22 22 1;
.print dc v(1,2) v(2,3) v(3);
.print dc i(vsupply);
.end;