*My own circuit with constant current source and 3 resistors in series

i1 1 0 dc 1.5e-3;
r1 1 2 4k;
r2 2 3 2k;
r3 3 0 5k;

.dc i1 1.5e-3 1.5e-3 1;
.print dc v(1,2) v(2,3) v(3);
.print dc v(1,0);
.end;